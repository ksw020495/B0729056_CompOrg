library verilog;
use verilog.vl_types.all;
entity b0729056_lab02 is
    port(
        X0              : in     vl_logic;
        X1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic;
        clk             : in     vl_logic;
        clean           : in     vl_logic;
        A0              : out    vl_logic;
        A1              : out    vl_logic;
        A2              : out    vl_logic;
        A3              : out    vl_logic;
        L               : out    vl_logic;
        A4u             : out    vl_logic
    );
end b0729056_lab02;
