library verilog;
use verilog.vl_types.all;
entity \7447\ is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        BIN             : in     vl_logic;
        LTN             : in     vl_logic;
        RBIN            : in     vl_logic;
        OG              : out    vl_logic;
        \OF\            : out    vl_logic;
        OE              : out    vl_logic;
        RBON            : out    vl_logic;
        OD              : out    vl_logic;
        OC              : out    vl_logic;
        OB              : out    vl_logic;
        OA              : out    vl_logic
    );
end \7447\;
