library verilog;
use verilog.vl_types.all;
entity lab05 is
    port(
        Count           : in     vl_logic;
        clk             : in     vl_logic;
        clean           : in     vl_logic;
        Q0A             : out    vl_logic;
        Q0B             : out    vl_logic;
        Q0C             : out    vl_logic;
        Q0D             : out    vl_logic;
        Q0E             : out    vl_logic;
        Q0F             : out    vl_logic;
        Q0G             : out    vl_logic;
        Q1A             : out    vl_logic;
        Q1B             : out    vl_logic;
        Q1C             : out    vl_logic;
        Q1D             : out    vl_logic;
        Q1E             : out    vl_logic;
        Q1F             : out    vl_logic;
        Q1G             : out    vl_logic;
        Q2A             : out    vl_logic;
        Q2B             : out    vl_logic;
        Q2C             : out    vl_logic;
        Q2D             : out    vl_logic;
        Q2E             : out    vl_logic;
        Q2F             : out    vl_logic;
        Q2G             : out    vl_logic;
        Q3A             : out    vl_logic;
        Q3B             : out    vl_logic;
        Q3C             : out    vl_logic;
        Q3D             : out    vl_logic;
        Q3E             : out    vl_logic;
        Q3F             : out    vl_logic;
        Q3G             : out    vl_logic
    );
end lab05;
